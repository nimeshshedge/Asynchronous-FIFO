module wptr_full (
 output reg wfull,
 output [4-1:0] waddr,
 output reg [4 :0] wptr,
 input [4 :0] wq2_rptr,
 input winc, wclk, wrst_n);
 
 reg [4:0] wbin;
 wire [4:0] wgraynext, wbinnext;
 
 // GRAYSTYLE2 pointer
 always @(posedge wclk or negedge wrst_n)
	if (!wrst_n) 
		{wbin, wptr} <= 0;
	else 
		{wbin, wptr} <= {wbinnext, wgraynext};
 
 // Memory write-address pointer (okay to use binary to address memory)
 assign waddr = wbin[4-1:0];
 assign wbinnext = wbin + (winc & ~wfull);
 assign wgraynext = (wbinnext>>1) ^ wbinnext;
 
 //------------------------------------------------------------------
 // Simplified version of the three necessary full-tests:
 // assign wfull_val=((wgnext[ADDRSIZE] !=wq2_rptr[ADDRSIZE] ) &&
 // (wgnext[ADDRSIZE-1] !=wq2_rptr[ADDRSIZE-1]) &&
 // (wgnext[ADDRSIZE-2:0]==wq2_rptr[ADDRSIZE-2:0]));
 //------------------------------------------------------------------

 assign wfull_val = (wgraynext=={~wq2_rptr[4:4-1], wq2_rptr[4-2:0]});
 always @(posedge wclk or negedge wrst_n)
	if (!wrst_n) 
		wfull <= 1'b0;
	else 
		wfull <= wfull_val;
		
endmodule